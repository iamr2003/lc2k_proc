module imem(
    input [31:0] pc, //I'll just assume it's an integer like everything else
    output [31:0] instr
);
// need to figure out how to load this properly
// functions similar to normal memory, just has no writing

endmodule
