module imem()
// need to figure out how to load this properly

endmodule
